module alu_datapath(clk, alu_data_a, alu_data_b, store_a, store_b, start_alu, finished, result, overflow)






module bit_parity(bit_a, bit_b, bit_parity_out)

input bit_a;
input bit_b;
input bit_borrow_in;

output bit_diff;
output bit_borrow_out;
module bit_subtractor(bit_a, bit_b, bit_borrow_in, bit_diff, bit_borrow_out)

input bit_a;
input bit_b;
input bit_borrow_in;

output bit_diff;
output bit_borrow_out;

module top();



endmodule